module Program_Counter
  
(
  input [63:0] PC_In,
  output reg [63:0] PC_Out,
  input clk,
  input reset
);


always @ (posedge reset or posedge clk)

begin
  
if (reset)
  assign PC_Out = 64'h0000000000000000;

else
  assign PC_Out = PC_In;
  
end

endmodule
